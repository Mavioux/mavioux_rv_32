module mavioux_rv_32 (
    
)