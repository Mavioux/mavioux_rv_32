module mavioux_rv_32 (
    
);

endmodule